module vdl 

struct C.SDL_Surface {}

pub struct Surface {
	ptr &C.SDL_Surface
}