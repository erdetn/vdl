module vdl 

struct C.SDL_Surface {}

pub fn Surface {
	ptr &C.SDL_Surface
}